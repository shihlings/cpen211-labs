module regfile(data_in,writenum,write,readnum,clk,data_out);
   input [15:0] data_in;
   input [2:0]	writenum, readnum;
   input	write, clk;
   output [15:0] data_out;
   // fill out the rest
endmodule
