module shifter(in,shift,sout);
   input [15:0] in;
   input [1:0]	shift;
   output [15:0] sout;
   // fill out the rest
endmodule
