module tb_lab3();
// hello
endmodule: tb_lab3
