module datapath;
   
endmodule // datapath
